`include "define.v"

module memory(
    input  wire        clk_i,
    input  wire [ 2:0] M_stat_i,
    input  wire [ 3:0] M_icode_i,
    input  wire [63:0] M_valE_i,
    input  wire [63:0] M_valA_i,
    input  wire [ 3:0] M_dstE_i,
    input  wire [ 3:0] M_dstM_i,

    output wire [ 2:0] m_stat_o,
    output wire [63:0] m_valM_o
);

wire        mem_read;
wire        mem_write;
wire        dmem_error;
wire [63:0] addr;

assign mem_read = (M_icode_i == `IMRMOVQ) | (M_icode_i == `IPOPQ) | (M_icode_i == `IRET);
assign mem_write = (M_icode_i == `IRMMOVQ) | (M_icode_i == `IPUSHQ) | (M_icode_i == `ICALL);
assign addr =  (M_icode_i == `IRMMOVQ || M_icode_i == `IMRMOVQ || 
            M_icode_i == `IPUSHQ || M_icode_i == `ICALL) ? M_valE_i : 
            (M_icode_i == `IPOPQ || M_icode_i == `IRET) ? M_valA_i : 64'b0;
assign m_stat_o = dmem_error ? `SADR : M_stat_i;
ram mem(
    .clk_i(clk_i),
    .addr_i(addr),
    .data_i(M_valA_i),
    .read_i(mem_read),
    .write_i(mem_write),
    .dmem_error_o(dmem_error),
    .data_o(m_valM_o)
);
endmodule

module ram (
    input  wire        clk_i,
    input  wire [63:0] addr_i,
    input  wire [63:0] data_i,
    input  wire        read_i,
    input  wire        write_i,

    output wire        dmem_error_o,
    output wire [63:0] data_o
);

parameter MAX_SIZE = 1024;
reg [7:0] mem[0:1023];

assign dmem_error_o = (addr_i >= MAX_SIZE) ? 1 : 0;

always @(posedge clk_i) begin
    if (write_i) { mem[addr_i + 7], mem[addr_i + 6], 
    mem[addr_i + 5], mem[addr_i + 4],
    mem[addr_i + 3], mem[addr_i + 2],
    mem[addr_i + 1], mem[addr_i] } <= data_i;
end

assign data_o = read_i ? { mem[addr_i + 7], mem[addr_i + 6], 
    mem[addr_i + 5], mem[addr_i + 4],
    mem[addr_i + 3], mem[addr_i + 2],
    mem[addr_i + 1], mem[addr_i] } : 64'b0;

initial begin
//                            | # Array of 4 elements
//0x018:                      | 	.align 8
//0x018: 0100000001000000     | array:	.quad 0x0000000100000001
    mem[24] = 8'h01;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h01;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
//0x020: 0100000001000000     | 	.quad 0x0000000100000001
    mem[32] = 8'h01;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h01;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
//0x028: 0100000001000000     | 	.quad 0x0000000100000001
    mem[40] = 8'h01;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h01;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
//0x030: 0100000001000000     | 	.quad 0x0000000100000001
    mem[48] = 8'h01;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h01;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
//0x038: 0100000001000000     | 	.quad 0x0000000100000001
    mem[56] = 8'h01;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h01;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
//0x040: 0100000001000000     | 	.quad 0x0000000100000001
    mem[64] = 8'h01;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h01;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
//0x048: 0100000001000000     | 	.quad 0x0000000100000001
    mem[72] = 8'h01;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h01;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
//0x050: 0100000001000000     | 	.quad 0x0000000100000001
    mem[80] = 8'h01;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h01;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
//0x058: 0100000001000000     | 	.quad 0x0000000100000001
    mem[88] = 8'h01;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h01;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
//0x060: 0100000001000000     | 	.quad 0x0000000100000001
    mem[96] = 8'h01;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h01;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
//0x068: 0100000001000000     | 	.quad 0x0000000100000001
    mem[104] = 8'h01;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h01;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
//0x070: 0100000001000000     | 	.quad 0x0000000100000001
    mem[112] = 8'h01;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h01;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
//0x078: 0100000001000000     | 	.quad 0x0000000100000001
    mem[120] = 8'h01;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h01;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
//0x080: 0100000001000000     | 	.quad 0x0000000100000001
    mem[128] = 8'h01;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h01;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
//0x088: 0100000001000000     | 	.quad 0x0000000100000001
    mem[136] = 8'h01;
    mem[137] = 8'h00;
    mem[138] = 8'h00;
    mem[139] = 8'h00;
    mem[140] = 8'h01;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
//0x090: 0100000001000000     | 	.quad 0x0000000100000001
    mem[144] = 8'h01;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'h00;
    mem[148] = 8'h01;
    mem[149] = 8'h00;
    mem[150] = 8'h00;
    mem[151] = 8'h00;
//0x098: 0100000001000000     | 	.quad 0x0000000100000001
    mem[152] = 8'h01;
    mem[153] = 8'h00;
    mem[154] = 8'h00;
    mem[155] = 8'h00;
    mem[156] = 8'h01;
    mem[157] = 8'h00;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
//0x0a0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[160] = 8'h01;
    mem[161] = 8'h00;
    mem[162] = 8'h00;
    mem[163] = 8'h00;
    mem[164] = 8'h01;
    mem[165] = 8'h00;
    mem[166] = 8'h00;
    mem[167] = 8'h00;
//0x0a8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[168] = 8'h01;
    mem[169] = 8'h00;
    mem[170] = 8'h00;
    mem[171] = 8'h00;
    mem[172] = 8'h01;
    mem[173] = 8'h00;
    mem[174] = 8'h00;
    mem[175] = 8'h00;
//0x0b0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[176] = 8'h01;
    mem[177] = 8'h00;
    mem[178] = 8'h00;
    mem[179] = 8'h00;
    mem[180] = 8'h01;
    mem[181] = 8'h00;
    mem[182] = 8'h00;
    mem[183] = 8'h00;
//0x0b8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[184] = 8'h01;
    mem[185] = 8'h00;
    mem[186] = 8'h00;
    mem[187] = 8'h00;
    mem[188] = 8'h01;
    mem[189] = 8'h00;
    mem[190] = 8'h00;
    mem[191] = 8'h00;
//0x0c0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[192] = 8'h01;
    mem[193] = 8'h00;
    mem[194] = 8'h00;
    mem[195] = 8'h00;
    mem[196] = 8'h01;
    mem[197] = 8'h00;
    mem[198] = 8'h00;
    mem[199] = 8'h00;
//0x0c8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[200] = 8'h01;
    mem[201] = 8'h00;
    mem[202] = 8'h00;
    mem[203] = 8'h00;
    mem[204] = 8'h01;
    mem[205] = 8'h00;
    mem[206] = 8'h00;
    mem[207] = 8'h00;
//0x0d0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[208] = 8'h01;
    mem[209] = 8'h00;
    mem[210] = 8'h00;
    mem[211] = 8'h00;
    mem[212] = 8'h01;
    mem[213] = 8'h00;
    mem[214] = 8'h00;
    mem[215] = 8'h00;
//0x0d8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[216] = 8'h01;
    mem[217] = 8'h00;
    mem[218] = 8'h00;
    mem[219] = 8'h00;
    mem[220] = 8'h01;
    mem[221] = 8'h00;
    mem[222] = 8'h00;
    mem[223] = 8'h00;
//0x0e0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[224] = 8'h01;
    mem[225] = 8'h00;
    mem[226] = 8'h00;
    mem[227] = 8'h00;
    mem[228] = 8'h01;
    mem[229] = 8'h00;
    mem[230] = 8'h00;
    mem[231] = 8'h00;
//0x0e8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[232] = 8'h01;
    mem[233] = 8'h00;
    mem[234] = 8'h00;
    mem[235] = 8'h00;
    mem[236] = 8'h01;
    mem[237] = 8'h00;
    mem[238] = 8'h00;
    mem[239] = 8'h00;
//0x0f0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[240] = 8'h01;
    mem[241] = 8'h00;
    mem[242] = 8'h00;
    mem[243] = 8'h00;
    mem[244] = 8'h01;
    mem[245] = 8'h00;
    mem[246] = 8'h00;
    mem[247] = 8'h00;
//0x0f8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[248] = 8'h01;
    mem[249] = 8'h00;
    mem[250] = 8'h00;
    mem[251] = 8'h00;
    mem[252] = 8'h01;
    mem[253] = 8'h00;
    mem[254] = 8'h00;
    mem[255] = 8'h00;
//0x100: 0100000001000000     | 	.quad 0x0000000100000001
    mem[256] = 8'h01;
    mem[257] = 8'h00;
    mem[258] = 8'h00;
    mem[259] = 8'h00;
    mem[260] = 8'h01;
    mem[261] = 8'h00;
    mem[262] = 8'h00;
    mem[263] = 8'h00;
//0x108: 0100000001000000     | 	.quad 0x0000000100000001
    mem[264] = 8'h01;
    mem[265] = 8'h00;
    mem[266] = 8'h00;
    mem[267] = 8'h00;
    mem[268] = 8'h01;
    mem[269] = 8'h00;
    mem[270] = 8'h00;
    mem[271] = 8'h00;
//0x110: 0100000001000000     | 	.quad 0x0000000100000001
    mem[272] = 8'h01;
    mem[273] = 8'h00;
    mem[274] = 8'h00;
    mem[275] = 8'h00;
    mem[276] = 8'h01;
    mem[277] = 8'h00;
    mem[278] = 8'h00;
    mem[279] = 8'h00;
//0x118: 0100000001000000     | 	.quad 0x0000000100000001
    mem[280] = 8'h01;
    mem[281] = 8'h00;
    mem[282] = 8'h00;
    mem[283] = 8'h00;
    mem[284] = 8'h01;
    mem[285] = 8'h00;
    mem[286] = 8'h00;
    mem[287] = 8'h00;
//0x120: 0100000001000000     | 	.quad 0x0000000100000001
    mem[288] = 8'h01;
    mem[289] = 8'h00;
    mem[290] = 8'h00;
    mem[291] = 8'h00;
    mem[292] = 8'h01;
    mem[293] = 8'h00;
    mem[294] = 8'h00;
    mem[295] = 8'h00;
//0x128: 0100000001000000     | 	.quad 0x0000000100000001
    mem[296] = 8'h01;
    mem[297] = 8'h00;
    mem[298] = 8'h00;
    mem[299] = 8'h00;
    mem[300] = 8'h01;
    mem[301] = 8'h00;
    mem[302] = 8'h00;
    mem[303] = 8'h00;
//0x130: 0100000001000000     | 	.quad 0x0000000100000001
    mem[304] = 8'h01;
    mem[305] = 8'h00;
    mem[306] = 8'h00;
    mem[307] = 8'h00;
    mem[308] = 8'h01;
    mem[309] = 8'h00;
    mem[310] = 8'h00;
    mem[311] = 8'h00;
//0x138: 0100000001000000     | 	.quad 0x0000000100000001
    mem[312] = 8'h01;
    mem[313] = 8'h00;
    mem[314] = 8'h00;
    mem[315] = 8'h00;
    mem[316] = 8'h01;
    mem[317] = 8'h00;
    mem[318] = 8'h00;
    mem[319] = 8'h00;
//0x140: 0100000001000000     | 	.quad 0x0000000100000001
    mem[320] = 8'h01;
    mem[321] = 8'h00;
    mem[322] = 8'h00;
    mem[323] = 8'h00;
    mem[324] = 8'h01;
    mem[325] = 8'h00;
    mem[326] = 8'h00;
    mem[327] = 8'h00;
//0x148: 0100000001000000     | 	.quad 0x0000000100000001
    mem[328] = 8'h01;
    mem[329] = 8'h00;
    mem[330] = 8'h00;
    mem[331] = 8'h00;
    mem[332] = 8'h01;
    mem[333] = 8'h00;
    mem[334] = 8'h00;
    mem[335] = 8'h00;
//0x150: 0100000001000000     | 	.quad 0x0000000100000001
    mem[336] = 8'h01;
    mem[337] = 8'h00;
    mem[338] = 8'h00;
    mem[339] = 8'h00;
    mem[340] = 8'h01;
    mem[341] = 8'h00;
    mem[342] = 8'h00;
    mem[343] = 8'h00;
//0x158: 0100000001000000     | 	.quad 0x0000000100000001
    mem[344] = 8'h01;
    mem[345] = 8'h00;
    mem[346] = 8'h00;
    mem[347] = 8'h00;
    mem[348] = 8'h01;
    mem[349] = 8'h00;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
//0x160: 0100000001000000     | 	.quad 0x0000000100000001
    mem[352] = 8'h01;
    mem[353] = 8'h00;
    mem[354] = 8'h00;
    mem[355] = 8'h00;
    mem[356] = 8'h01;
    mem[357] = 8'h00;
    mem[358] = 8'h00;
    mem[359] = 8'h00;
//0x168: 0100000001000000     | 	.quad 0x0000000100000001
    mem[360] = 8'h01;
    mem[361] = 8'h00;
    mem[362] = 8'h00;
    mem[363] = 8'h00;
    mem[364] = 8'h01;
    mem[365] = 8'h00;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
//0x170: 0100000001000000     | 	.quad 0x0000000100000001
    mem[368] = 8'h01;
    mem[369] = 8'h00;
    mem[370] = 8'h00;
    mem[371] = 8'h00;
    mem[372] = 8'h01;
    mem[373] = 8'h00;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
//0x178: 0100000001000000     | 	.quad 0x0000000100000001
    mem[376] = 8'h01;
    mem[377] = 8'h00;
    mem[378] = 8'h00;
    mem[379] = 8'h00;
    mem[380] = 8'h01;
    mem[381] = 8'h00;
    mem[382] = 8'h00;
    mem[383] = 8'h00;
//0x180: 0100000001000000     | 	.quad 0x0000000100000001
    mem[384] = 8'h01;
    mem[385] = 8'h00;
    mem[386] = 8'h00;
    mem[387] = 8'h00;
    mem[388] = 8'h01;
    mem[389] = 8'h00;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
//0x188: 0100000001000000     | 	.quad 0x0000000100000001
    mem[392] = 8'h01;
    mem[393] = 8'h00;
    mem[394] = 8'h00;
    mem[395] = 8'h00;
    mem[396] = 8'h01;
    mem[397] = 8'h00;
    mem[398] = 8'h00;
    mem[399] = 8'h00;
//0x190: 0100000001000000     | 	.quad 0x0000000100000001
    mem[400] = 8'h01;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h01;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
//0x198: 0100000001000000     | 	.quad 0x0000000100000001
    mem[408] = 8'h01;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h01;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
//0x1a0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[416] = 8'h01;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h01;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
//0x1a8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[424] = 8'h01;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h01;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
//0x1b0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[432] = 8'h01;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h01;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
//0x1b8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[440] = 8'h01;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h01;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
//0x1c0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[448] = 8'h01;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h01;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
//0x1c8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[456] = 8'h01;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h01;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
//0x1d0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[464] = 8'h01;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h01;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
//0x1d8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[472] = 8'h01;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h01;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
//0x1e0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[480] = 8'h01;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h01;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
//0x1e8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[488] = 8'h01;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h01;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
//0x1f0: 0100000001000000     | 	.quad 0x0000000100000001
    mem[496] = 8'h01;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h01;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
//0x1f8: 0100000001000000     | 	.quad 0x0000000100000001
    mem[504] = 8'h01;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h01;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
//0x200: 0100000001000000     | 	.quad 0x0000000100000001
    mem[512] = 8'h01;
    mem[513] = 8'h00;
    mem[514] = 8'h00;
    mem[515] = 8'h00;
    mem[516] = 8'h01;
    mem[517] = 8'h00;
    mem[518] = 8'h00;
    mem[519] = 8'h00;
//0x208: 0100000001000000     | 	.quad 0x0000000100000001
    mem[520] = 8'h01;
    mem[521] = 8'h00;
    mem[522] = 8'h00;
    mem[523] = 8'h00;
    mem[524] = 8'h01;
    mem[525] = 8'h00;
    mem[526] = 8'h00;
    mem[527] = 8'h00;
//0x210: 0100000001000000     | 	.quad 0x0000000100000001
    mem[528] = 8'h01;
    mem[529] = 8'h00;
    mem[530] = 8'h00;
    mem[531] = 8'h00;
    mem[532] = 8'h01;
    mem[533] = 8'h00;
    mem[534] = 8'h00;
    mem[535] = 8'h00;
//                            | 
end
endmodule